// softproc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module softproc (
		input  wire        clk_clk,                                   //                       clk.clk
		input  wire        master_template_0_control_fixed_location,  // master_template_0_control.fixed_location
		input  wire [31:0] master_template_0_control_write_base,      //                          .write_base
		input  wire [31:0] master_template_0_control_write_length,    //                          .write_length
		input  wire        master_template_0_control_go,              //                          .go
		output wire        master_template_0_control_done,            //                          .done
		input  wire        master_template_0_user_write_buffer,       //    master_template_0_user.write_buffer
		input  wire [31:0] master_template_0_user_buffer_input_data,  //                          .buffer_input_data
		output wire        master_template_0_user_buffer_full,        //                          .buffer_full
		input  wire        master_template_1_control_fixed_location,  // master_template_1_control.fixed_location
		input  wire [31:0] master_template_1_control_read_base,       //                          .read_base
		input  wire [31:0] master_template_1_control_read_length,     //                          .read_length
		input  wire        master_template_1_control_go,              //                          .go
		output wire        master_template_1_control_done,            //                          .done
		output wire        master_template_1_control_early_done,      //                          .early_done
		input  wire        master_template_1_user_read_buffer,        //    master_template_1_user.read_buffer
		output wire [31:0] master_template_1_user_buffer_output_data, //                          .buffer_output_data
		output wire        master_template_1_user_data_available,     //                          .data_available
		output wire        sdram_clock_clk,                           //               sdram_clock.clk
		output wire [12:0] sdram_wire_addr,                           //                sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                          .ba
		output wire        sdram_wire_cas_n,                          //                          .cas_n
		output wire        sdram_wire_cke,                            //                          .cke
		output wire        sdram_wire_cs_n,                           //                          .cs_n
		inout  wire [31:0] sdram_wire_dq,                             //                          .dq
		output wire [3:0]  sdram_wire_dqm,                            //                          .dqm
		output wire        sdram_wire_ras_n,                          //                          .ras_n
		output wire        sdram_wire_we_n                            //                          .we_n
	);

	wire         sys_sdram_pll_0_sys_clk_clk;                                 // sys_sdram_pll_0:sys_clk_clk -> [irq_mapper:clk, jtag_uart_0:clk, master_template_0:clk, master_template_1:clk, mm_interconnect_0:sys_sdram_pll_0_sys_clk_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_003:reset_in1]
	wire         master_template_0_avalon_master_waitrequest;                 // mm_interconnect_0:master_template_0_avalon_master_waitrequest -> master_template_0:master_waitrequest
	wire  [31:0] master_template_0_avalon_master_address;                     // master_template_0:master_address -> mm_interconnect_0:master_template_0_avalon_master_address
	wire   [3:0] master_template_0_avalon_master_byteenable;                  // master_template_0:master_byteenable -> mm_interconnect_0:master_template_0_avalon_master_byteenable
	wire         master_template_0_avalon_master_write;                       // master_template_0:master_write -> mm_interconnect_0:master_template_0_avalon_master_write
	wire  [31:0] master_template_0_avalon_master_writedata;                   // master_template_0:master_writedata -> mm_interconnect_0:master_template_0_avalon_master_writedata
	wire  [31:0] master_template_1_avalon_master_readdata;                    // mm_interconnect_0:master_template_1_avalon_master_readdata -> master_template_1:master_readdata
	wire         master_template_1_avalon_master_waitrequest;                 // mm_interconnect_0:master_template_1_avalon_master_waitrequest -> master_template_1:master_waitrequest
	wire  [31:0] master_template_1_avalon_master_address;                     // master_template_1:master_address -> mm_interconnect_0:master_template_1_avalon_master_address
	wire         master_template_1_avalon_master_read;                        // master_template_1:master_read -> mm_interconnect_0:master_template_1_avalon_master_read
	wire   [3:0] master_template_1_avalon_master_byteenable;                  // master_template_1:master_byteenable -> mm_interconnect_0:master_template_1_avalon_master_byteenable
	wire         master_template_1_avalon_master_readdatavalid;               // mm_interconnect_0:master_template_1_avalon_master_readdatavalid -> master_template_1:master_readdatavalid
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;      // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;        // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;     // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;         // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;            // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [3:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;      // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;   // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;           // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [31:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;       // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, master_template_0:reset, master_template_1:reset, mm_interconnect_0:master_template_0_clock_reset_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> onchip_memory2_0:reset_req
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> sys_sdram_pll_0:ref_reset_reset

	softproc_jtag_uart_0 jtag_uart_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                                 //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	custom_master #(
		.MASTER_DIRECTION    (1),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) master_template_0 (
		.clk                     (sys_sdram_pll_0_sys_clk_clk),                 //       clock_reset.clk
		.reset                   (rst_controller_001_reset_out_reset),          // clock_reset_reset.reset
		.master_address          (master_template_0_avalon_master_address),     //     avalon_master.address
		.master_write            (master_template_0_avalon_master_write),       //                  .write
		.master_byteenable       (master_template_0_avalon_master_byteenable),  //                  .byteenable
		.master_writedata        (master_template_0_avalon_master_writedata),   //                  .writedata
		.master_waitrequest      (master_template_0_avalon_master_waitrequest), //                  .waitrequest
		.control_fixed_location  (master_template_0_control_fixed_location),    //           control.export
		.control_write_base      (master_template_0_control_write_base),        //                  .export
		.control_write_length    (master_template_0_control_write_length),      //                  .export
		.control_go              (master_template_0_control_go),                //                  .export
		.control_done            (master_template_0_control_done),              //                  .export
		.user_write_buffer       (master_template_0_user_write_buffer),         //              user.export
		.user_buffer_input_data  (master_template_0_user_buffer_input_data),    //                  .export
		.user_buffer_full        (master_template_0_user_buffer_full),          //                  .export
		.master_read             (),                                            //       (terminated)
		.master_readdata         (32'b00000000000000000000000000000000),        //       (terminated)
		.master_readdatavalid    (1'b0),                                        //       (terminated)
		.master_burstcount       (),                                            //       (terminated)
		.control_read_base       (32'b00000000000000000000000000000000),        //       (terminated)
		.control_read_length     (32'b00000000000000000000000000000000),        //       (terminated)
		.control_early_done      (),                                            //       (terminated)
		.user_read_buffer        (1'b0),                                        //       (terminated)
		.user_buffer_output_data (),                                            //       (terminated)
		.user_data_available     ()                                             //       (terminated)
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (0),
		.MAXIMUM_BURST_COUNT (2),
		.BURST_COUNT_WIDTH   (2),
		.FIFO_DEPTH          (32),
		.FIFO_DEPTH_LOG2     (5),
		.MEMORY_BASED_FIFO   (1)
	) master_template_1 (
		.clk                     (sys_sdram_pll_0_sys_clk_clk),                   //       clock_reset.clk
		.reset                   (rst_controller_001_reset_out_reset),            // clock_reset_reset.reset
		.master_address          (master_template_1_avalon_master_address),       //     avalon_master.address
		.master_read             (master_template_1_avalon_master_read),          //                  .read
		.master_byteenable       (master_template_1_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (master_template_1_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (master_template_1_avalon_master_readdatavalid), //                  .readdatavalid
		.master_waitrequest      (master_template_1_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (master_template_1_control_fixed_location),      //           control.export
		.control_read_base       (master_template_1_control_read_base),           //                  .export
		.control_read_length     (master_template_1_control_read_length),         //                  .export
		.control_go              (master_template_1_control_go),                  //                  .export
		.control_done            (master_template_1_control_done),                //                  .export
		.control_early_done      (master_template_1_control_early_done),          //                  .export
		.user_read_buffer        (master_template_1_user_read_buffer),            //              user.export
		.user_buffer_output_data (master_template_1_user_buffer_output_data),     //                  .export
		.user_data_available     (master_template_1_user_data_available),         //                  .export
		.master_write            (),                                              //       (terminated)
		.master_writedata        (),                                              //       (terminated)
		.master_burstcount       (),                                              //       (terminated)
		.control_write_base      (32'b00000000000000000000000000000000),          //       (terminated)
		.control_write_length    (32'b00000000000000000000000000000000),          //       (terminated)
		.user_write_buffer       (1'b0),                                          //       (terminated)
		.user_buffer_input_data  (32'b00000000000000000000000000000000),          //       (terminated)
		.user_buffer_full        ()                                               //       (terminated)
	);

	softproc_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (sys_sdram_pll_0_sys_clk_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                           //  wire.export
		.zs_ba          (sdram_wire_ba),                                             //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                          //      .export
		.zs_cke         (sdram_wire_cke),                                            //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                           //      .export
		.zs_dq          (sdram_wire_dq),                                             //      .export
		.zs_dqm         (sdram_wire_dqm),                                            //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                          //      .export
		.zs_we_n        (sdram_wire_we_n)                                            //      .export
	);

	softproc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sys_sdram_pll_0_sys_clk_clk),                                //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	softproc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sys_sdram_pll_0_sys_clk_clk),                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	softproc_sys_sdram_pll_0 sys_sdram_pll_0 (
		.ref_clk_clk        (clk_clk),                            //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_sdram_pll_0_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clock_clk),                    //    sdram_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	softproc_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_0_sys_clk_clk                                     (sys_sdram_pll_0_sys_clk_clk),                                 //                                   sys_sdram_pll_0_sys_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                              //                   jtag_uart_0_reset_reset_bridge_in_reset.reset
		.master_template_0_clock_reset_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // master_template_0_clock_reset_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                          //             onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.master_template_0_avalon_master_address                         (master_template_0_avalon_master_address),                     //                           master_template_0_avalon_master.address
		.master_template_0_avalon_master_waitrequest                     (master_template_0_avalon_master_waitrequest),                 //                                                          .waitrequest
		.master_template_0_avalon_master_byteenable                      (master_template_0_avalon_master_byteenable),                  //                                                          .byteenable
		.master_template_0_avalon_master_write                           (master_template_0_avalon_master_write),                       //                                                          .write
		.master_template_0_avalon_master_writedata                       (master_template_0_avalon_master_writedata),                   //                                                          .writedata
		.master_template_1_avalon_master_address                         (master_template_1_avalon_master_address),                     //                           master_template_1_avalon_master.address
		.master_template_1_avalon_master_waitrequest                     (master_template_1_avalon_master_waitrequest),                 //                                                          .waitrequest
		.master_template_1_avalon_master_byteenable                      (master_template_1_avalon_master_byteenable),                  //                                                          .byteenable
		.master_template_1_avalon_master_read                            (master_template_1_avalon_master_read),                        //                                                          .read
		.master_template_1_avalon_master_readdata                        (master_template_1_avalon_master_readdata),                    //                                                          .readdata
		.master_template_1_avalon_master_readdatavalid                   (master_template_1_avalon_master_readdatavalid),               //                                                          .readdatavalid
		.nios2_gen2_0_data_master_address                                (nios2_gen2_0_data_master_address),                            //                                  nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                            (nios2_gen2_0_data_master_waitrequest),                        //                                                          .waitrequest
		.nios2_gen2_0_data_master_byteenable                             (nios2_gen2_0_data_master_byteenable),                         //                                                          .byteenable
		.nios2_gen2_0_data_master_read                                   (nios2_gen2_0_data_master_read),                               //                                                          .read
		.nios2_gen2_0_data_master_readdata                               (nios2_gen2_0_data_master_readdata),                           //                                                          .readdata
		.nios2_gen2_0_data_master_write                                  (nios2_gen2_0_data_master_write),                              //                                                          .write
		.nios2_gen2_0_data_master_writedata                              (nios2_gen2_0_data_master_writedata),                          //                                                          .writedata
		.nios2_gen2_0_data_master_debugaccess                            (nios2_gen2_0_data_master_debugaccess),                        //                                                          .debugaccess
		.nios2_gen2_0_instruction_master_address                         (nios2_gen2_0_instruction_master_address),                     //                           nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                     (nios2_gen2_0_instruction_master_waitrequest),                 //                                                          .waitrequest
		.nios2_gen2_0_instruction_master_read                            (nios2_gen2_0_instruction_master_read),                        //                                                          .read
		.nios2_gen2_0_instruction_master_readdata                        (nios2_gen2_0_instruction_master_readdata),                    //                                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_address                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                             jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                          .write
		.jtag_uart_0_avalon_jtag_slave_read                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                          .read
		.jtag_uart_0_avalon_jtag_slave_readdata                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                          .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                          .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                          .chipselect
		.new_sdram_controller_0_s1_address                               (mm_interconnect_0_new_sdram_controller_0_s1_address),         //                                 new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                                 (mm_interconnect_0_new_sdram_controller_0_s1_write),           //                                                          .write
		.new_sdram_controller_0_s1_read                                  (mm_interconnect_0_new_sdram_controller_0_s1_read),            //                                                          .read
		.new_sdram_controller_0_s1_readdata                              (mm_interconnect_0_new_sdram_controller_0_s1_readdata),        //                                                          .readdata
		.new_sdram_controller_0_s1_writedata                             (mm_interconnect_0_new_sdram_controller_0_s1_writedata),       //                                                          .writedata
		.new_sdram_controller_0_s1_byteenable                            (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),      //                                                          .byteenable
		.new_sdram_controller_0_s1_readdatavalid                         (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),   //                                                          .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                           (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),     //                                                          .waitrequest
		.new_sdram_controller_0_s1_chipselect                            (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),      //                                                          .chipselect
		.nios2_gen2_0_debug_mem_slave_address                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //                              nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                                          .write
		.nios2_gen2_0_debug_mem_slave_read                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                                          .read
		.nios2_gen2_0_debug_mem_slave_readdata                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                                          .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                                          .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                                          .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                                          .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                                          .debugaccess
		.onchip_memory2_0_s1_address                                     (mm_interconnect_0_onchip_memory2_0_s1_address),               //                                       onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                       (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                                          .write
		.onchip_memory2_0_s1_readdata                                    (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                                          .readdata
		.onchip_memory2_0_s1_writedata                                   (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                                          .writedata
		.onchip_memory2_0_s1_byteenable                                  (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                                          .byteenable
		.onchip_memory2_0_s1_chipselect                                  (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                                          .chipselect
		.onchip_memory2_0_s1_clken                                       (mm_interconnect_0_onchip_memory2_0_s1_clken)                  //                                                          .clken
	);

	softproc_irq_mapper irq_mapper (
		.clk           (sys_sdram_pll_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (sys_sdram_pll_0_sys_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
